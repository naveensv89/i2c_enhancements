module test();

initial
  $display("Hello World!");
  
endmodule
